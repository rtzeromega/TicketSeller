module FOUR_in(led,a,b,c,d);
	output led;
	input a,b,c,d;
	reg led,tmp1,tmp2;
	
	always @(a or b or c or d)
	begin
	 tmp1=a&b;
	 tmp2=c&d;
	 led=~(tmp1|tmp2);
	end
endmodule
